`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   12:21:08 04/04/2023
// Design Name:   sync_3bit_upcounter
// Module Name:   /home/jay711/VERILOG_CODES/COUNTERS/sync_3bit_upcounter_tb.v
// Project Name:  COUNTERS
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: sync_3bit_upcounter
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module sync_3bit_upcounter_tb;

	// Inputs
	reg clk;
	reg rst;

	// Outputs
	wire [2:0] q;

	// Instantiate the Unit Under Test (UUT)
	sync_3bit_upcounter uut (
		.clk(clk), 
		.rst(rst), 
		.q(q)
	);

initial begin
		clk = 1; rst = 1;
		#10; clk=1; rst=0;
	end
	
	always
	forever #5 clk=~clk;
	
	initial begin
	$monitor("time=%g clk=%b rst=%b count=%b",$time,clk,rst,q);
	#2000 $finish;
	end
      
endmodule

